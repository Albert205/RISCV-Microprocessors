import Opcode_pkg::*;

class OpCode_class;
    randc OpCode_t OpCode;
endclass
