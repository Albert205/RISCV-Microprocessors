package ALUControl_pkg;
    typedef enum bit[2:0] {ADD = 3'd0, SUB = 3'd1, AND = 3'd2, OR = 3'd3, SLT = 3'd5} ALUControl_t;

endpackage : ALUControl_pkg